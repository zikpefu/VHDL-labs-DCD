LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY comparator IS
port(A: IN STD_LOGIC_VECTOR(15 downto 0);
B: IN STD_LOGIC_VECTOR(15 downto 0);
O: OUT STD_LOGIC);
END comparator;

ARCHITECTURE behavior OF comparator  IS
begin
end behavior;